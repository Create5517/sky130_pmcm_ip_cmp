** sch_path: /home/kali/Desktop/Chipalooza_April2024_Comparator/cace/input_offset.sch
**.subckt input_offset
Vavdd avdd VSUB DC 3.3
Rout vout VSUB 100000000.0 m=1
Cout vout VSUB 1e-13 m=1
Vdvdd dvdd VSUB DC 1.8
?
?
Vavss avss VSUB DC 0
Vdvss dvss VSUB DC 0
RSUB VSUB GND 0.01 m=1
Iibias VSUB ibias DC 1e-06
XDUT hsyt_0 hsyt_1 avdd vinp avss vinn dvdd dvss vout ibias ena Chipalooza_April2024_Comparator
?
?
VVcm inx VSUB DC {Vcm}
**** begin user architecture code

* CACE gensim simulation file inputOffset_1
* Generated by CACE gensim, Efabless Corporation (c) 2023
* Find the current through the amplifier under condition of static input

.include ./netlist/schematic/Chipalooza_April2024_Comparator.spice


.lib /usr/local/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice ss

.option TEMP=27
* Flag unsafe operating conditions (exceeds models' specified limits)
.option warn=1
.option savecurrents
.option save all



.control
** Find zero crossing for positive input differential, zero crossing for negative
** input differential, then compute the average
tran [{risetime} * 2 / 1000] [{risetime} * 2]
meas tran vhigh FIND V(inp) WHEN V(out) = [{Vvdd} / 2] CROSS=1
meas tran vlow FIND V(inp) WHEN V(out) = [{Vvdd} / 2] CROSS=2
let vrise = $&vhigh - {Vcm}
let vfall = $&vlow - {Vcm}

let voffset = 0.5 * ($&vrise + $&vfall)
let vhyst = $&vrise - $&vfall

echo $&voffset $&vhyst > ngspice/inputOffset_1.data
*set wr_singlescale
*wrdata ngspice/inputOffset_1.data V(out) V(inp) V(inm)

write ngspice/input_offset.raw

quit
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
