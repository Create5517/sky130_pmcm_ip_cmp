** sch_path: /home/kali/Desktop/Chipalooza_April2024_Comparator/cace/input_offset.sch
**.subckt input_offset
Vavdd avdd VSUB DC {Vavdd}
Rout vout VSUB {Rout} m=1
Cout vout VSUB {Cout} m=1
Vdvdd dvdd VSUB DC {Vdvdd}
?
?
Vavss avss VSUB DC {Vavss}
Vdvss dvss VSUB DC {Vdvss}
RSUB VSUB GND 0.01 m=1
Iibias VSUB ibias DC {ibias}
XDUT hsyt_0 hsyt_1 avdd vinp avss vinn dvdd dvss vout ibias ena Chipalooza_April2024_Comparator
?
?
VVcm inx VSUB DC {Vcm}
**** begin user architecture code

* CACE gensim simulation file {filename}_{N}
* Generated by CACE gensim, Efabless Corporation (c) 2023
* Find the current through the amplifier under condition of static input

.include {DUT_path}

.lib {PDK_ROOT}/{PDK}/libs.tech/combined/sky130.lib.spice {corner}

.option TEMP={temperature}
* Flag unsafe operating conditions (exceeds models' specified limits)
.option warn=1
.option savecurrents
.option save all



.control
** Find zero crossing for positive input differential, zero crossing for negative
** input differential, then compute the average
tran [{risetime} * 2 / 1000] [{risetime} * 2]
meas tran vhigh FIND V(inp) WHEN V(out) = [{Vvdd} / 2] CROSS=1
meas tran vlow FIND V(inp) WHEN V(out) = [{Vvdd} / 2] CROSS=2
let vrise = $&vhigh - {Vcm}
let vfall = $&vlow - {Vcm}

let voffset = 0.5 * ($&vrise + $&vfall)
let vhyst = $&vrise - $&vfall

echo $&voffset $&vhyst > {simpath}/{filename}_{N}.data
*set wr_singlescale
*wrdata {simpath}/{filename}_{N}.data V(out) V(inp) V(inm)

write ngspice/input_offset.raw

quit
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
