** sch_path: /home/kali/Desktop/ZacMayGit/OLD8_sky130_pmcm_ip_cmp/Chipalooza_April2024_Comparator/xschem/Chipalooza_April2024_Comparator.sch
.subckt Chipalooza_April2024_Comparator vinp vinn hyst0 hyst1 avdd avss dvdd dvss vout ena ibias
*.PININFO vinp:I vinn:I hyst0:I hyst1:I avdd:I avss:I dvdd:I dvss:I vout:O ena:I ibias:I
C1 avss 0 2p m=1
XEN avssi ena avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=4 nf=1 m=4
XHS_IB1 net3 ibias avssi avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 m=2
XOS_P2 vout SumOutBar dvdd dvdd sky130_fd_pr__pfet_01v8 L=1 W=2 nf=1 m=2
XOS_N2 vout SumOutBar avssi dvss sky130_fd_pr__nfet_01v8 L=1 W=2 nf=1 m=2
XSC_P1 SourceBias2 SourceBias2 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 m=2
XSC_P2 N1 SourceBias2 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 m=2
XSC_P3 N2 SourceBias2 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 m=2
XSC_p5 SumOut Bias1 N2 avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 m=2
XSC_P4 Sum Bias1 N1 avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 m=2
XSC_N2 SumOut Bias2 P2 avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=2
XSC_N1 Sum Bias2 P1 avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=2
XSC_N4 P2 Sum avssi avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=2
XSC_N3 P1 Sum avssi avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=2
XIS_PIN2 P2 vinn psource_input avdd sky130_fd_pr__pfet_g5v0d10v5 L=4 W=32 nf=1 m=2
XIS_PIN1 P1 vinp psource_input avdd sky130_fd_pr__pfet_g5v0d10v5 L=4 W=32 nf=1 m=2
XIS_PMIR3X psource_input net4 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=12 nf=1 m=4
XIS_PMIR1X net4 net4 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=8 nf=1 m=2
XIS_PSWITCH nbias_tail net9 psource_input avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=8 nf=1 m=2
XIS_NIN1 N1 vinp SourceBias0 avss sky130_fd_pr__nfet_g5v0d10v5 L=4 W=16 nf=1 m=2
XIS_NIN2 N2 vinn SourceBias0 avss sky130_fd_pr__nfet_g5v0d10v5 L=4 W=16 nf=1 m=2
XIS_NMIR3X SourceBias0 nbias_tail avssi avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=12 nf=1 m=4
XIS_NMIR1X nbias_tail nbias_tail avssi avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=12 nf=1 m=2
XIS_NSWITCH net4 Bias5 SourceBias0 avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=4 nf=1 m=2
XCM_SB1 SourceBias1 ibias avssi avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=3 nf=1 m=2
XIS_PIREF1 SourceBias1 SourceBias1 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=12 nf=1 m=4
XIS_PIREF2 psource_input SourceBias1 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=12 nf=1 m=4
XCM_SB2 SourceBias2 ibias avssi avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=6 nf=1 m=2
XCM_SB3 SourceBias3 ibias avssi avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 m=2
XCM_BIAS1 Bias1 ibias avssi avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=3 nf=1 m=2
XCM_SB5 SourceBias5 ibias avssi avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=3 nf=1 m=2
XCM_SB6 SourceBias6 ibias avssi avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=3 nf=1 m=2
XCM_SB7 SourceBias7 ibias avssi avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=3 nf=1 m=2
XCM_BIAS5 Bias5 ibias avssi avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=3 nf=1 m=2
XB2_N3 M55Source M55Drain avssi avss sky130_fd_pr__nfet_g5v0d10v5 L=1.5 W=6 nf=1 m=2
XB2_N1 M55Drain Bias2 M55Source avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=9 nf=1 m=2
XB2_N2 Bias2 Bias2 avssi avss sky130_fd_pr__nfet_g5v0d10v5 L=2 W=0.5 nf=1 m=1
XB1_P1 net5 net6 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=2 W=20 nf=1 m=2
XB1_P2 net6 net6 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=2 W=10 nf=1 m=2
XB1_P5 SourceBias4 SourceBias4 net6 avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=10 nf=1 m=2
XB1_P4 avssi SourceBias4 net5 avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1 nf=1 m=2
XB1_P3 Bias1 Bias1 net5 avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=5 nf=1 m=2
XB5_P1 net7 net8 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=2 W=20 nf=1 m=2
XB5_P2 net8 net8 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=2 W=20 nf=1 m=2
XB5_P5 SourceBias7 SourceBias7 net8 avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=10 nf=1 m=2
XB5_P4 avssi SourceBias7 net7 avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1 nf=1 m=2
XB5_P3 Bias5 Bias5 net7 avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=5 nf=1 m=2
XB2_P1 SourceBias5 SourceBias5 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=12 nf=1 m=4
XB2_P2 M55Drain SourceBias5 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=12 nf=1 m=4
XB2_P4 SourceBias6 SourceBias6 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=12 nf=1 m=4
XB2_P3 Bias2 SourceBias6 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=12 nf=1 m=4
XCM_SB0 SourceBias0 ibias avssi avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=3 nf=1 m=2
XHS_N1 N1 SumOut net1 avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=2
XHS_N2 N2 SumOutBar net1 avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=2
XIB_N1 ibias ibias avssi avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=3 nf=1 m=2
XIB_N2 avdd ibias avssi avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=3 nf=1 m=2
XIS_PSWITCH_B3 net9 net9 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=5 W=3 nf=1 m=1
XIS_PSWTICH_B1 avdd Bias4 SourceBias3 avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=4 nf=1 m=2
XIS_PSWITCH_B2 net9 Bias5 SourceBias3 avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=4 nf=1 m=2
XB4_P1 net10 net11 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=2 W=20 nf=1 m=2
XB4_P2 net11 net11 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=2 W=10 nf=1 m=2
XB4_P5 SourceBias10 SourceBias10 net11 avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=10 nf=1 m=2
XM1 net2 ibias avssi avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 m=2
XHS_H0 net1 hyst0 net2 avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 m=2
XHS_H1 net1 hyst1 net3 avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=2
XCM_BIAS4 Bias4 ibias avssi avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=3 nf=1 m=2
XCM_SB10 SourceBias10 ibias avssi avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=3 nf=1 m=2
XCM_SB4 SourceBias4 ibias avssi avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=3 nf=1 m=2
XB4_P4 avssi SourceBias10 net10 avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1 nf=1 m=2
XB4_P3 Bias4 Bias4 net10 avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=5 nf=1 m=2
XM29 SumOutBar SumOut dvdd dvdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 m=2
XM30 SumOutBar SumOut avssi dvss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=2
.ends
.end
