** sch_path: /home/kali/Desktop/Chipalooza_April2024_Comparator/cace/powerConsumption.sch
**.subckt powerConsumption
Vavdd avdd VSUB DC {Vavdd}
Rout vout VSUB {Rout} m=1
Cout vout VSUB {Cout} m=1
Vdvdd dvdd VSUB DC {Vdvdd}
Vvcm vinn VSUB DC {Vvcm}
Vena ena VSUB DC {ena}
Vhyst0 hyst0 VSUB DC 1.8
Vavss avss VSUB DC {Vavss}
Vdvss dvss VSUB DC {Vdvss}
RSUB VSUB GND 0.01 m=1
Iibias VSUB ibias DC {ibias}
VVdiff vinp vinn DC {Vdiff}
XDUT hyst0 hyst1 avdd vinp avss vinn dvdd dvss vout ibias ena Chipalooza_April2024_Comparator
Vhyst1 hyst1 VSUB DC 1.8
**** begin user architecture code

.control
op

set wr_singlescale
wrdata {simpath}/{filename}_{N}.data -I(Vdvdd)
write ngspice/powerConsumption.raw

quit

.endc



* CACE gensim simulation file {filename}_{N}
* Generated by CACE gensim, Efabless Corporation (c) 2023
* Find the current through the amplifier under condition of static input

.include {DUT_path}

.lib {PDK_ROOT}/{PDK}/libs.tech/combined/sky130.lib.spice {corner}

.option TEMP={temperature}
* Flag unsafe operating conditions (exceeds models' specified limits)
.option warn=1
.option savecurrents
.option save all


**** end user architecture code
**.ends
.GLOBAL GND
.end
