** sch_path: /home/kali/Desktop/Chipalooza_April2024_Comparator/cace/cmrr.sch
**.subckt cmrr
Vavdd avdd VSUB DC {Vavdd}
Rout vout VSUB {Rout} m=1
Cout vout VSUB {Cout} m=1
Vdvdd dvdd VSUB DC {Vdvdd}
?
?
Vavss avss VSUB DC {Vavss}
Vdvss dvss VSUB DC {Vdvss}
RSUB VSUB GND 0.01 m=1
Iibias VSUB ibias DC {ibias}
XDUT hsyt_0 hsyt_1 avdd vinp avss vinn dvdd dvss vout ibias ena Chipalooza_April2024_Comparator
?
?
?
**** begin user architecture code

.control
** CMRR is defined as the change in input offset vs. change in common-mode voltage.
tran [{risetime} * 2 / 100] [{risetime} * 4]
meas tran vhigh1 FIND V(vinp) WHEN V(vout) = [{Vavdd} / 2] CROSS=1
meas tran vlow1 FIND V(vinp) WHEN V(vout) = [{Vavdd} / 2] CROSS=2
meas tran vhigh2 FIND V(vinp) WHEN V(vout) = [{Vavdd} / 2] CROSS=3
meas tran vlow2 FIND V(vinp) WHEN V(vout) = [{Vavdd} / 2] CROSS=4

let voffset1 = 0.5 * ($&vhigh1 + $&vlow1) - {Vcm|minimum}
let voffset2 = 0.5 * ($&vhigh2 + $&vlow2) - {Vcm|maximum}

let cmrr = ($&voffset1 - $&voffset2) / ({Vcm|maximum} - {Vcm|minimum})
let cmrrdb = 20 * log(abs($&cmrr))

echo $&cmrrdb > {simpath}/{filename}_{N}.data

write ngspice/cmrr.raw

quit
.endc



* CACE gensim simulation file {filename}_{N}
* Generated by CACE gensim, Efabless Corporation (c) 2023
* Find the power supply rejection ratio of the amplifier

.include {DUT_path}

.lib {PDK_ROOT}/{PDK}/libs.tech/combined/sky130.lib.spice {corner}

.option TEMP={temperature}
* Flag unsafe operating conditions (exceeds models' specified limits)
.option warn=1
.option savecurrents
.option save all


**** end user architecture code
**.ends
.GLOBAL GND
.end
