** sch_path: /home/kali/Desktop/Chipalooza_April2024_Comparator/cace/powerConsumption.sch
.subckt powerConsumption

Vavdd avdd VSUB DC {Vavdd}
Rout vout VSUB {Rout} m=1
Cout vout VSUB {Cout} m=1
Vdvdd dvdd VSUB DC {Vdvdd}
Vvcm vinn VSUB DC {Vvcm}
?
?
Vavss avss VSUB DC {Vavss}
Vdvss dvss VSUB DC {Vdvss}
RSUB VSUB GND 0.01 m=1
Iibias VSUB ibias DC {ibias}
VVdiff vinp vinn DC {Vdiff}
x1 hsyt_0 hsyt_1 avdd vinp avss vinn dvdd dvss vout ibias ena Chipalooza_April2024_Comparator
**** begin user architecture code

.control
option savecurrents
op
set wr_singlescale
wrdata {simpath}/{filename}_{N}.data -I(Vdvdd)
write ngspice/powerConsumption.raw
quit
.endc



* CACE gensim simulation file {filename}_{N}
* Generated by CACE gensim, Efabless Corporation (c) 2023
* Find the current through the amplifier under condition of static input

.include {DUT_path}

.lib {PDK_ROOT}/{PDK}/libs.tech/combined/sky130.lib.spice {corner}

.option TEMP={temperature}
* Flag unsafe operating conditions (exceeds models' specified limits)
.option warn=1
.option savecurrents
.option save all


**** end user architecture code
.ends

* expanding   symbol:  /home/kali/Desktop/Chipalooza_April2024_Comparator/xschem/Chipalooza_April2024_Comparator.sym # of pins=11
** sym_path: /home/kali/Desktop/Chipalooza_April2024_Comparator/xschem/Chipalooza_April2024_Comparator.sym
** sch_path: /home/kali/Desktop/Chipalooza_April2024_Comparator/xschem/Chipalooza_April2024_Comparator.sch
.subckt Chipalooza_April2024_Comparator vhyst_0 vhyst_1 avdd vinp avss vinn dvdd dvss vout ibias ena
*.PININFO vinp:I vinn:I vhyst_0:I vhyst_1:I avdd:I avss:I dvdd:I dvss:I vout:O ena:I ibias:I
XM1 ibias ibias net3 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 net2 ibias net3 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 net1 vinp net2 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 net5 vinn net2 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 I_hyst I_hyst net3 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 net1 vout net4 dvss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 net4 I_hyst net3 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM8 net5 net6 net4 dvss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM9 net6 ibias net3 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM11 net1 net1 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM12 net5 net1 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM15 net6 net5 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM13 ibias vhyst_0 net8 dvss sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
C38 avss 0 2p m=1
XM24 net3 ena avss avss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM16 ibias vhyst_1 net7 dvss sky130_fd_pr__nfet_01v8 L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM19 net7 vhyst_bias I_hyst dvss sky130_fd_pr__nfet_01v8 L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM18 net8 vhyst_bias I_hyst dvss sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM10 vout net6 net3 avss sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM14 vout net6 dvdd dvdd sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
V1 vhyst_bias GND 1.2
.ends

.GLOBAL GND
.end
