** sch_path: /home/kali/Desktop/Chipalooza_April2024_Comparator/cace/frequencyBandwidth.sch
**.subckt frequencyBandwidth
Vavdd avdd VSUB DC {Vavdd}
Rout vout VSUB {Rout} m=1
Cout vout VSUB {Cout} m=1
Vdvdd dvdd VSUB DC {Vdvdd}
?
?
?
Vavss avss VSUB DC {Vavss}
Vdvss dvss VSUB DC {Vdvss}
RSUB VSUB GND 0.01 m=1
Iibias VSUB ibias DC {ibias}
XDUT vhyst_0 vhyst_1 avdd vinp avss vinn dvdd dvss vout ibias ena Chipalooza_April2024_Comparator
VVpos vinp inx DC 1.65 AC 1.65
VVneg inx vinn DC -1.65
VVcm inx VSUB DC {Vcm}
**** begin user architecture code

.control

ac dec 20 1 1e12
plot v(vout)
plot v(dvdd)
plot v(avdd)

meas ac peak MAX vmag(vout) FROM=2 TO=1.5GHz
let f3db = peak/sqrt(2)
meas ac f1 when vmag(vout)=f3db RISE=1
meas ac f2 when vmag(vout)=f3db FALL=1

let f3 = $&f2
echo $&f3 > {simpath}/{filename}_{N}.data

write ngspice/frequencyBandwidth.raw

.endc



* CACE gensim simulation file {filename}_{N}
* Generated by CACE gensim, Efabless Corporation (c) 2023
* Find the current through the amplifier under condition of static input

.include {DUT_path}

.lib {PDK_ROOT}/{PDK}/libs.tech/combined/sky130.lib.spice {corner}

.option TEMP={temperature}
* Flag unsafe operating conditions (exceeds models' specified limits)
.option warn=1
.option savecurrents
.option save all


**** end user architecture code
**.ends
.GLOBAL GND
.end
